// megafunction wizard: %LPM_DECODE%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_decode 

// ============================================================
// File Name: lpm_decode1.v
// Megafunction Name(s):
// 			lpm_decode
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 222 10/21/2009 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module lpm_decode1 (
	data,
	eq00,
	eq01,
	eq02,
	eq03,
	eq04,
	eq05,
	eq06,
	eq07,
	eq08,
	eq09,
	eq0a,
	eq0b,
	eq0c,
	eq0d,
	eq0e,
	eq0f);

	input	[3:0]  data;
	output	  eq00;
	output	  eq01;
	output	  eq02;
	output	  eq03;
	output	  eq04;
	output	  eq05;
	output	  eq06;
	output	  eq07;
	output	  eq08;
	output	  eq09;
	output	  eq0a;
	output	  eq0b;
	output	  eq0c;
	output	  eq0d;
	output	  eq0e;
	output	  eq0f;

	wire [15:0] sub_wire0;
	wire [4:4] sub_wire16 = sub_wire0[4:4];
	wire [14:14] sub_wire15 = sub_wire0[14:14];
	wire [3:3] sub_wire14 = sub_wire0[3:3];
	wire [13:13] sub_wire13 = sub_wire0[13:13];
	wire [2:2] sub_wire12 = sub_wire0[2:2];
	wire [12:12] sub_wire11 = sub_wire0[12:12];
	wire [1:1] sub_wire10 = sub_wire0[1:1];
	wire [11:11] sub_wire9 = sub_wire0[11:11];
	wire [0:0] sub_wire8 = sub_wire0[0:0];
	wire [10:10] sub_wire7 = sub_wire0[10:10];
	wire [9:9] sub_wire6 = sub_wire0[9:9];
	wire [8:8] sub_wire5 = sub_wire0[8:8];
	wire [7:7] sub_wire4 = sub_wire0[7:7];
	wire [6:6] sub_wire3 = sub_wire0[6:6];
	wire [5:5] sub_wire2 = sub_wire0[5:5];
	wire [15:15] sub_wire1 = sub_wire0[15:15];
	wire  eq0f = sub_wire1;
	wire  eq05 = sub_wire2;
	wire  eq06 = sub_wire3;
	wire  eq07 = sub_wire4;
	wire  eq08 = sub_wire5;
	wire  eq09 = sub_wire6;
	wire  eq0a = sub_wire7;
	wire  eq00 = sub_wire8;
	wire  eq0b = sub_wire9;
	wire  eq01 = sub_wire10;
	wire  eq0c = sub_wire11;
	wire  eq02 = sub_wire12;
	wire  eq0d = sub_wire13;
	wire  eq03 = sub_wire14;
	wire  eq0e = sub_wire15;
	wire  eq04 = sub_wire16;

	lpm_decode	lpm_decode_component (
				.data (data),
				.eq (sub_wire0)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock (),
				.enable ()
				// synopsys translate_on
				);
	defparam
		lpm_decode_component.lpm_decodes = 16,
		lpm_decode_component.lpm_type = "LPM_DECODE",
		lpm_decode_component.lpm_width = 4;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: BaseDec NUMERIC "0"
// Retrieval info: PRIVATE: EnableInput NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
// Retrieval info: PRIVATE: Latency NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: eq0 NUMERIC "1"
// Retrieval info: PRIVATE: eq1 NUMERIC "1"
// Retrieval info: PRIVATE: eq10 NUMERIC "1"
// Retrieval info: PRIVATE: eq11 NUMERIC "1"
// Retrieval info: PRIVATE: eq12 NUMERIC "1"
// Retrieval info: PRIVATE: eq13 NUMERIC "1"
// Retrieval info: PRIVATE: eq14 NUMERIC "1"
// Retrieval info: PRIVATE: eq15 NUMERIC "1"
// Retrieval info: PRIVATE: eq2 NUMERIC "1"
// Retrieval info: PRIVATE: eq3 NUMERIC "1"
// Retrieval info: PRIVATE: eq4 NUMERIC "1"
// Retrieval info: PRIVATE: eq5 NUMERIC "1"
// Retrieval info: PRIVATE: eq6 NUMERIC "1"
// Retrieval info: PRIVATE: eq7 NUMERIC "1"
// Retrieval info: PRIVATE: eq8 NUMERIC "1"
// Retrieval info: PRIVATE: eq9 NUMERIC "1"
// Retrieval info: PRIVATE: nBit NUMERIC "4"
// Retrieval info: CONSTANT: LPM_DECODES NUMERIC "16"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DECODE"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "4"
// Retrieval info: USED_PORT: @eq 0 0 LPM_DECODES 0 OUTPUT NODEFVAL @eq[LPM_DECODES-1..0]
// Retrieval info: USED_PORT: data 0 0 4 0 INPUT NODEFVAL data[3..0]
// Retrieval info: USED_PORT: eq00 0 0 0 0 OUTPUT NODEFVAL eq00
// Retrieval info: USED_PORT: eq01 0 0 0 0 OUTPUT NODEFVAL eq01
// Retrieval info: USED_PORT: eq02 0 0 0 0 OUTPUT NODEFVAL eq02
// Retrieval info: USED_PORT: eq03 0 0 0 0 OUTPUT NODEFVAL eq03
// Retrieval info: USED_PORT: eq04 0 0 0 0 OUTPUT NODEFVAL eq04
// Retrieval info: USED_PORT: eq05 0 0 0 0 OUTPUT NODEFVAL eq05
// Retrieval info: USED_PORT: eq06 0 0 0 0 OUTPUT NODEFVAL eq06
// Retrieval info: USED_PORT: eq07 0 0 0 0 OUTPUT NODEFVAL eq07
// Retrieval info: USED_PORT: eq08 0 0 0 0 OUTPUT NODEFVAL eq08
// Retrieval info: USED_PORT: eq09 0 0 0 0 OUTPUT NODEFVAL eq09
// Retrieval info: USED_PORT: eq0A 0 0 0 0 OUTPUT NODEFVAL eq0A
// Retrieval info: USED_PORT: eq0B 0 0 0 0 OUTPUT NODEFVAL eq0B
// Retrieval info: USED_PORT: eq0C 0 0 0 0 OUTPUT NODEFVAL eq0C
// Retrieval info: USED_PORT: eq0D 0 0 0 0 OUTPUT NODEFVAL eq0D
// Retrieval info: USED_PORT: eq0E 0 0 0 0 OUTPUT NODEFVAL eq0E
// Retrieval info: USED_PORT: eq0F 0 0 0 0 OUTPUT NODEFVAL eq0F
// Retrieval info: CONNECT: @data 0 0 4 0 data 0 0 4 0
// Retrieval info: CONNECT: eq00 0 0 0 0 @eq 0 0 1 0
// Retrieval info: CONNECT: eq01 0 0 0 0 @eq 0 0 1 1
// Retrieval info: CONNECT: eq02 0 0 0 0 @eq 0 0 1 2
// Retrieval info: CONNECT: eq03 0 0 0 0 @eq 0 0 1 3
// Retrieval info: CONNECT: eq04 0 0 0 0 @eq 0 0 1 4
// Retrieval info: CONNECT: eq05 0 0 0 0 @eq 0 0 1 5
// Retrieval info: CONNECT: eq06 0 0 0 0 @eq 0 0 1 6
// Retrieval info: CONNECT: eq07 0 0 0 0 @eq 0 0 1 7
// Retrieval info: CONNECT: eq08 0 0 0 0 @eq 0 0 1 8
// Retrieval info: CONNECT: eq09 0 0 0 0 @eq 0 0 1 9
// Retrieval info: CONNECT: eq0A 0 0 0 0 @eq 0 0 1 10
// Retrieval info: CONNECT: eq0B 0 0 0 0 @eq 0 0 1 11
// Retrieval info: CONNECT: eq0C 0 0 0 0 @eq 0 0 1 12
// Retrieval info: CONNECT: eq0D 0 0 0 0 @eq 0 0 1 13
// Retrieval info: CONNECT: eq0E 0 0 0 0 @eq 0 0 1 14
// Retrieval info: CONNECT: eq0F 0 0 0 0 @eq 0 0 1 15
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode1.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode1.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode1.cmp TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode1.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode1_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode1_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
